magic
tech sky130A
magscale 1 2
timestamp 1698610993
<< metal3 >>
rect -4492 6332 -120 6360
rect -4492 2308 -204 6332
rect -140 2308 -120 6332
rect -4492 2280 -120 2308
rect 120 6332 4492 6360
rect 120 2308 4408 6332
rect 4472 2308 4492 6332
rect 120 2280 4492 2308
rect -4492 2012 -120 2040
rect -4492 -2012 -204 2012
rect -140 -2012 -120 2012
rect -4492 -2040 -120 -2012
rect 120 2012 4492 2040
rect 120 -2012 4408 2012
rect 4472 -2012 4492 2012
rect 120 -2040 4492 -2012
rect -4492 -2308 -120 -2280
rect -4492 -6332 -204 -2308
rect -140 -6332 -120 -2308
rect -4492 -6360 -120 -6332
rect 120 -2308 4492 -2280
rect 120 -6332 4408 -2308
rect 4472 -6332 4492 -2308
rect 120 -6360 4492 -6332
<< via3 >>
rect -204 2308 -140 6332
rect 4408 2308 4472 6332
rect -204 -2012 -140 2012
rect 4408 -2012 4472 2012
rect -204 -6332 -140 -2308
rect 4408 -6332 4472 -2308
<< mimcap >>
rect -4452 6280 -452 6320
rect -4452 2360 -4412 6280
rect -492 2360 -452 6280
rect -4452 2320 -452 2360
rect 160 6280 4160 6320
rect 160 2360 200 6280
rect 4120 2360 4160 6280
rect 160 2320 4160 2360
rect -4452 1960 -452 2000
rect -4452 -1960 -4412 1960
rect -492 -1960 -452 1960
rect -4452 -2000 -452 -1960
rect 160 1960 4160 2000
rect 160 -1960 200 1960
rect 4120 -1960 4160 1960
rect 160 -2000 4160 -1960
rect -4452 -2360 -452 -2320
rect -4452 -6280 -4412 -2360
rect -492 -6280 -452 -2360
rect -4452 -6320 -452 -6280
rect 160 -2360 4160 -2320
rect 160 -6280 200 -2360
rect 4120 -6280 4160 -2360
rect 160 -6320 4160 -6280
<< mimcapcontact >>
rect -4412 2360 -492 6280
rect 200 2360 4120 6280
rect -4412 -1960 -492 1960
rect 200 -1960 4120 1960
rect -4412 -6280 -492 -2360
rect 200 -6280 4120 -2360
<< metal4 >>
rect -2504 6281 -2400 6480
rect -224 6332 -120 6480
rect -4413 6280 -491 6281
rect -4413 2360 -4412 6280
rect -492 2360 -491 6280
rect -4413 2359 -491 2360
rect -2504 1961 -2400 2359
rect -224 2308 -204 6332
rect -140 2308 -120 6332
rect 2108 6281 2212 6480
rect 4388 6332 4492 6480
rect 199 6280 4121 6281
rect 199 2360 200 6280
rect 4120 2360 4121 6280
rect 199 2359 4121 2360
rect -224 2012 -120 2308
rect -4413 1960 -491 1961
rect -4413 -1960 -4412 1960
rect -492 -1960 -491 1960
rect -4413 -1961 -491 -1960
rect -2504 -2359 -2400 -1961
rect -224 -2012 -204 2012
rect -140 -2012 -120 2012
rect 2108 1961 2212 2359
rect 4388 2308 4408 6332
rect 4472 2308 4492 6332
rect 4388 2012 4492 2308
rect 199 1960 4121 1961
rect 199 -1960 200 1960
rect 4120 -1960 4121 1960
rect 199 -1961 4121 -1960
rect -224 -2308 -120 -2012
rect -4413 -2360 -491 -2359
rect -4413 -6280 -4412 -2360
rect -492 -6280 -491 -2360
rect -4413 -6281 -491 -6280
rect -2504 -6480 -2400 -6281
rect -224 -6332 -204 -2308
rect -140 -6332 -120 -2308
rect 2108 -2359 2212 -1961
rect 4388 -2012 4408 2012
rect 4472 -2012 4492 2012
rect 4388 -2308 4492 -2012
rect 199 -2360 4121 -2359
rect 199 -6280 200 -2360
rect 4120 -6280 4121 -2360
rect 199 -6281 4121 -6280
rect -224 -6480 -120 -6332
rect 2108 -6480 2212 -6281
rect 4388 -6332 4408 -2308
rect 4472 -6332 4492 -2308
rect 4388 -6480 4492 -6332
<< properties >>
string FIXED_BBOX 120 2280 4200 6360
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

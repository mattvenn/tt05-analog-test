magic
tech sky130A
magscale 1 2
timestamp 1698599621
<< metal3 >>
rect -5492 7832 -120 7860
rect -5492 2808 -204 7832
rect -140 2808 -120 7832
rect -5492 2780 -120 2808
rect 120 7832 5492 7860
rect 120 2808 5408 7832
rect 5472 2808 5492 7832
rect 120 2780 5492 2808
rect -5492 2512 -120 2540
rect -5492 -2512 -204 2512
rect -140 -2512 -120 2512
rect -5492 -2540 -120 -2512
rect 120 2512 5492 2540
rect 120 -2512 5408 2512
rect 5472 -2512 5492 2512
rect 120 -2540 5492 -2512
rect -5492 -2808 -120 -2780
rect -5492 -7832 -204 -2808
rect -140 -7832 -120 -2808
rect -5492 -7860 -120 -7832
rect 120 -2808 5492 -2780
rect 120 -7832 5408 -2808
rect 5472 -7832 5492 -2808
rect 120 -7860 5492 -7832
<< via3 >>
rect -204 2808 -140 7832
rect 5408 2808 5472 7832
rect -204 -2512 -140 2512
rect 5408 -2512 5472 2512
rect -204 -7832 -140 -2808
rect 5408 -7832 5472 -2808
<< mimcap >>
rect -5452 7780 -452 7820
rect -5452 2860 -5412 7780
rect -492 2860 -452 7780
rect -5452 2820 -452 2860
rect 160 7780 5160 7820
rect 160 2860 200 7780
rect 5120 2860 5160 7780
rect 160 2820 5160 2860
rect -5452 2460 -452 2500
rect -5452 -2460 -5412 2460
rect -492 -2460 -452 2460
rect -5452 -2500 -452 -2460
rect 160 2460 5160 2500
rect 160 -2460 200 2460
rect 5120 -2460 5160 2460
rect 160 -2500 5160 -2460
rect -5452 -2860 -452 -2820
rect -5452 -7780 -5412 -2860
rect -492 -7780 -452 -2860
rect -5452 -7820 -452 -7780
rect 160 -2860 5160 -2820
rect 160 -7780 200 -2860
rect 5120 -7780 5160 -2860
rect 160 -7820 5160 -7780
<< mimcapcontact >>
rect -5412 2860 -492 7780
rect 200 2860 5120 7780
rect -5412 -2460 -492 2460
rect 200 -2460 5120 2460
rect -5412 -7780 -492 -2860
rect 200 -7780 5120 -2860
<< metal4 >>
rect -3004 7781 -2900 7980
rect -224 7832 -120 7980
rect -5413 7780 -491 7781
rect -5413 2860 -5412 7780
rect -492 2860 -491 7780
rect -5413 2859 -491 2860
rect -3004 2461 -2900 2859
rect -224 2808 -204 7832
rect -140 2808 -120 7832
rect 2608 7781 2712 7980
rect 5388 7832 5492 7980
rect 199 7780 5121 7781
rect 199 2860 200 7780
rect 5120 2860 5121 7780
rect 199 2859 5121 2860
rect -224 2512 -120 2808
rect -5413 2460 -491 2461
rect -5413 -2460 -5412 2460
rect -492 -2460 -491 2460
rect -5413 -2461 -491 -2460
rect -3004 -2859 -2900 -2461
rect -224 -2512 -204 2512
rect -140 -2512 -120 2512
rect 2608 2461 2712 2859
rect 5388 2808 5408 7832
rect 5472 2808 5492 7832
rect 5388 2512 5492 2808
rect 199 2460 5121 2461
rect 199 -2460 200 2460
rect 5120 -2460 5121 2460
rect 199 -2461 5121 -2460
rect -224 -2808 -120 -2512
rect -5413 -2860 -491 -2859
rect -5413 -7780 -5412 -2860
rect -492 -7780 -491 -2860
rect -5413 -7781 -491 -7780
rect -3004 -7980 -2900 -7781
rect -224 -7832 -204 -2808
rect -140 -7832 -120 -2808
rect 2608 -2859 2712 -2461
rect 5388 -2512 5408 2512
rect 5472 -2512 5492 2512
rect 5388 -2808 5492 -2512
rect 199 -2860 5121 -2859
rect 199 -7780 200 -2860
rect 5120 -7780 5121 -2860
rect 199 -7781 5121 -7780
rect -224 -7980 -120 -7832
rect 2608 -7980 2712 -7781
rect 5388 -7832 5408 -2808
rect 5472 -7832 5492 -2808
rect 5388 -7980 5492 -7832
<< properties >>
string FIXED_BBOX 120 2780 5200 7860
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25 l 25 val 1.269k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

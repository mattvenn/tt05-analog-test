VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_matt_divider_test
  CLASS BLOCK ;
  FOREIGN tt_um_matt_divider_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 157.320 BY 111.520 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.630 110.520 134.930 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 76.670 110.520 76.970 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 73.910 110.520 74.210 111.520 ;
        RECT 76.670 110.520 76.970 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 71.150 110.520 71.450 111.520 ;
        RECT 73.910 110.520 74.210 111.520 ;
        RECT 76.670 110.520 76.970 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 68.390 110.520 68.690 111.520 ;
        RECT 71.150 110.520 71.450 111.520 ;
        RECT 73.910 110.520 74.210 111.520 ;
        RECT 76.670 110.520 76.970 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 65.630 110.520 65.930 111.520 ;
        RECT 68.390 110.520 68.690 111.520 ;
        RECT 71.150 110.520 71.450 111.520 ;
        RECT 73.910 110.520 74.210 111.520 ;
        RECT 76.670 110.520 76.970 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END uo_out[7]
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 65.630 110.520 65.930 111.520 ;
        RECT 68.390 110.520 68.690 111.520 ;
        RECT 71.150 110.520 71.450 111.520 ;
        RECT 73.910 110.520 74.210 111.520 ;
        RECT 76.670 110.520 76.970 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
        RECT 38.360 2.990 63.950 106.180 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
        RECT 24.230 110.520 24.530 111.520 ;
        RECT 26.990 110.520 27.290 111.520 ;
        RECT 29.750 110.520 30.050 111.520 ;
        RECT 32.510 110.520 32.810 111.520 ;
        RECT 35.270 110.520 35.570 111.520 ;
        RECT 38.030 110.520 38.330 111.520 ;
        RECT 40.790 110.520 41.090 111.520 ;
        RECT 43.550 110.520 43.850 111.520 ;
        RECT 46.310 110.520 46.610 111.520 ;
        RECT 49.070 110.520 49.370 111.520 ;
        RECT 51.830 110.520 52.130 111.520 ;
        RECT 54.590 110.520 54.890 111.520 ;
        RECT 57.350 110.520 57.650 111.520 ;
        RECT 60.110 110.520 60.410 111.520 ;
        RECT 62.870 110.520 63.170 111.520 ;
        RECT 65.630 110.520 65.930 111.520 ;
        RECT 68.390 110.520 68.690 111.520 ;
        RECT 71.150 110.520 71.450 111.520 ;
        RECT 73.910 110.520 74.210 111.520 ;
        RECT 76.670 110.520 76.970 111.520 ;
        RECT 79.430 110.520 79.730 111.520 ;
        RECT 82.190 110.520 82.490 111.520 ;
        RECT 84.950 110.520 85.250 111.520 ;
        RECT 87.710 110.520 88.010 111.520 ;
        RECT 90.470 110.520 90.770 111.520 ;
        RECT 93.230 110.520 93.530 111.520 ;
        RECT 95.990 110.520 96.290 111.520 ;
        RECT 98.750 110.520 99.050 111.520 ;
        RECT 101.510 110.520 101.810 111.520 ;
        RECT 104.270 110.520 104.570 111.520 ;
        RECT 107.030 110.520 107.330 111.520 ;
        RECT 109.790 110.520 110.090 111.520 ;
        RECT 112.550 110.520 112.850 111.520 ;
        RECT 115.310 110.520 115.610 111.520 ;
        RECT 118.070 110.520 118.370 111.520 ;
        RECT 120.830 110.520 121.130 111.520 ;
        RECT 123.590 110.520 123.890 111.520 ;
        RECT 126.350 110.520 126.650 111.520 ;
        RECT 129.110 110.520 129.410 111.520 ;
        RECT 131.870 110.520 132.170 111.520 ;
        RECT 134.630 110.520 134.930 111.520 ;
        RECT 137.390 110.520 137.690 111.520 ;
        RECT 38.360 2.990 63.950 106.180 ;
        RECT 113.050 4.240 138.640 107.430 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 76.080 89.700 81.960 94.550 ;
      LAYER met1 ;
        RECT 71.170 89.530 89.630 99.790 ;
      LAYER met2 ;
        RECT 70.700 97.440 90.320 100.290 ;
      LAYER met3 ;
        RECT 70.850 97.370 90.240 100.520 ;
      LAYER met4 ;
        RECT 63.950 110.120 65.230 110.790 ;
        RECT 66.330 110.120 67.990 110.790 ;
        RECT 69.090 110.120 70.750 110.790 ;
        RECT 71.850 110.120 73.510 110.790 ;
        RECT 74.610 110.120 76.270 110.790 ;
        RECT 77.370 110.120 79.030 110.790 ;
        RECT 80.130 110.120 81.790 110.790 ;
        RECT 82.890 110.120 84.550 110.790 ;
        RECT 85.650 110.120 87.310 110.790 ;
        RECT 88.410 110.120 90.070 110.790 ;
        RECT 91.170 110.120 92.830 110.790 ;
        RECT 93.930 110.120 95.590 110.790 ;
        RECT 96.690 110.120 98.350 110.790 ;
        RECT 99.450 110.120 101.110 110.790 ;
        RECT 102.210 110.120 103.870 110.790 ;
        RECT 104.970 110.120 106.630 110.790 ;
        RECT 107.730 110.120 109.390 110.790 ;
        RECT 110.490 110.120 112.150 110.790 ;
        RECT 63.950 107.830 113.050 110.120 ;
        RECT 63.950 106.580 112.650 107.830 ;
        RECT 64.350 94.840 112.650 106.580 ;
  END
END tt_um_matt_divider_test
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1698571942
<< metal1 >>
rect -990 1914 -638 1988
rect -990 1638 -960 1914
rect -668 1638 -638 1914
rect -990 1582 -638 1638
rect -168 1924 184 1988
rect -168 1666 -128 1924
rect 124 1716 184 1924
rect 1564 1960 1916 2004
rect 124 1666 134 1716
rect -168 1582 134 1666
rect 1564 1702 1604 1960
rect 1856 1702 1916 1960
rect 1564 1598 1916 1702
rect 2316 1940 2668 1978
rect 2316 1682 2376 1940
rect 2628 1682 2668 1940
rect -924 -74 -654 1582
rect -152 1276 128 1582
rect 1614 1478 1856 1598
rect 2316 1572 2668 1682
rect -148 834 -28 1276
rect 1614 1080 1866 1478
rect 2374 1286 2652 1572
rect -152 422 10 834
rect 66 792 228 836
rect 1648 792 1850 1080
rect 66 622 1854 792
rect 66 424 228 622
rect 1648 582 1850 622
rect -450 -74 -86 66
rect -924 -306 -86 -74
rect -924 -358 -654 -306
rect -450 -350 -86 -306
rect -38 -140 124 76
rect 182 -60 546 78
rect 2374 -60 2644 1286
rect -38 -336 128 -140
rect -12 -492 128 -336
rect 182 -338 2644 -60
rect 416 -348 2644 -338
rect 2374 -374 2644 -348
rect -12 -522 1208 -492
rect -12 -656 1010 -522
rect 1164 -656 1208 -522
rect -12 -686 1208 -656
rect -12 -698 128 -686
<< via1 >>
rect -960 1638 -668 1914
rect -128 1666 124 1924
rect 1604 1702 1856 1960
rect 2376 1682 2628 1940
rect 1010 -656 1164 -522
<< metal2 >>
rect -1084 1914 -554 2018
rect -1084 1638 -960 1914
rect -668 1638 -554 1914
rect -1084 1538 -554 1638
rect -222 1924 308 2052
rect -222 1666 -128 1924
rect 124 1666 308 1924
rect -222 1572 308 1666
rect 664 1806 1194 2062
rect 1548 1960 2078 2102
rect 664 1582 1200 1806
rect 1548 1702 1604 1960
rect 1856 1702 2078 1960
rect 1548 1622 2078 1702
rect 2310 1940 2840 2108
rect 2310 1682 2376 1940
rect 2628 1682 2840 1940
rect 2310 1628 2840 1682
rect 958 -522 1200 1582
rect 958 -656 1010 -522
rect 1164 -656 1200 -522
rect 958 -698 1200 -656
use sky130_fd_pr__res_generic_po_D4RDDB  sky130_fd_pr__res_generic_po_D4RDDB_0
timestamp 1698571942
transform 1 0 39 0 1 251
box -195 -595 195 595
<< labels >>
rlabel metal2 -1084 1538 -960 2018 1 1
rlabel metal2 -222 1924 308 2052 1 2
rlabel metal2 664 1944 1194 2062 1 3
rlabel metal2 1548 1960 2078 2102 1 4
rlabel metal2 2310 1940 2840 2108 1 5
<< end >>

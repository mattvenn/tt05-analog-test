magic
tech sky130A
magscale 1 2
timestamp 1698571942
<< poly >>
rect -195 579 -129 595
rect -195 545 -179 579
rect -145 545 -129 579
rect -195 165 -129 545
rect -195 -545 -129 -165
rect -195 -579 -179 -545
rect -145 -579 -129 -545
rect -195 -595 -129 -579
rect -87 579 -21 595
rect -87 545 -71 579
rect -37 545 -21 579
rect -87 165 -21 545
rect -87 -545 -21 -165
rect -87 -579 -71 -545
rect -37 -579 -21 -545
rect -87 -595 -21 -579
rect 21 579 87 595
rect 21 545 37 579
rect 71 545 87 579
rect 21 165 87 545
rect 21 -545 87 -165
rect 21 -579 37 -545
rect 71 -579 87 -545
rect 21 -595 87 -579
rect 129 579 195 595
rect 129 545 145 579
rect 179 545 195 579
rect 129 165 195 545
rect 129 -545 195 -165
rect 129 -579 145 -545
rect 179 -579 195 -545
rect 129 -595 195 -579
<< polycont >>
rect -179 545 -145 579
rect -179 -579 -145 -545
rect -71 545 -37 579
rect -71 -579 -37 -545
rect 37 545 71 579
rect 37 -579 71 -545
rect 145 545 179 579
rect 145 -579 179 -545
<< npolyres >>
rect -195 -165 -129 165
rect -87 -165 -21 165
rect 21 -165 87 165
rect 129 -165 195 165
<< locali >>
rect -195 545 -179 579
rect -145 545 -129 579
rect -87 545 -71 579
rect -37 545 -21 579
rect 21 545 37 579
rect 71 545 87 579
rect 129 545 145 579
rect 179 545 195 579
rect -195 -579 -179 -545
rect -145 -579 -129 -545
rect -87 -579 -71 -545
rect -37 -579 -21 -545
rect 21 -579 37 -545
rect 71 -579 87 -545
rect 129 -579 145 -545
rect 179 -579 195 -545
<< viali >>
rect -179 545 -145 579
rect -71 545 -37 579
rect 37 545 71 579
rect 145 545 179 579
rect -179 182 -145 545
rect -71 182 -37 545
rect 37 182 71 545
rect 145 182 179 545
rect -179 -545 -145 -182
rect -71 -545 -37 -182
rect 37 -545 71 -182
rect 145 -545 179 -182
rect -179 -579 -145 -545
rect -71 -579 -37 -545
rect 37 -579 71 -545
rect 145 -579 179 -545
<< metal1 >>
rect -185 579 -139 591
rect -185 182 -179 579
rect -145 182 -139 579
rect -185 170 -139 182
rect -77 579 -31 591
rect -77 182 -71 579
rect -37 182 -31 579
rect -77 170 -31 182
rect 31 579 77 591
rect 31 182 37 579
rect 71 182 77 579
rect 31 170 77 182
rect 139 579 185 591
rect 139 182 145 579
rect 179 182 185 579
rect 139 170 185 182
rect -185 -182 -139 -170
rect -185 -579 -179 -182
rect -145 -579 -139 -182
rect -185 -591 -139 -579
rect -77 -182 -31 -170
rect -77 -579 -71 -182
rect -37 -579 -31 -182
rect -77 -591 -31 -579
rect 31 -182 77 -170
rect 31 -579 37 -182
rect 71 -579 77 -182
rect 31 -591 77 -579
rect 139 -182 185 -170
rect 139 -579 145 -182
rect 179 -579 185 -182
rect 139 -591 185 -579
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 1.650 m 1 nx 4 wmin 0.330 lmin 1.650 rho 48.2 val 241.0 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1698509327
<< metal1 >>
rect -990 1914 -638 1988
rect -990 1638 -960 1914
rect -668 1638 -638 1914
rect -990 1582 -638 1638
rect -168 1924 184 1988
rect -168 1666 -128 1924
rect 124 1716 184 1924
rect 722 1944 1074 2008
rect 722 1836 796 1944
rect 490 1752 796 1836
rect 124 1666 218 1716
rect -168 1582 218 1666
rect -900 336 -752 1582
rect 134 964 218 1582
rect 466 1686 796 1752
rect 1048 1686 1074 1944
rect 466 1612 1074 1686
rect 466 1054 618 1612
rect 722 1602 1074 1612
rect 1564 1960 1916 2004
rect 1564 1702 1604 1960
rect 1856 1702 1916 1960
rect 1564 1598 1916 1702
rect 2316 1940 2668 1978
rect 2316 1682 2376 1940
rect 2628 1682 2668 1940
rect 1614 1326 1856 1598
rect 2316 1572 2668 1682
rect 916 1206 1856 1326
rect 906 1132 1856 1206
rect -88 564 426 964
rect 486 356 570 1054
rect 906 964 1024 1132
rect 1614 1128 1856 1132
rect 634 534 1228 964
rect -906 322 -178 336
rect -906 14 178 322
rect -360 -44 178 14
rect 278 -30 826 356
rect 1024 322 1618 350
rect 2440 322 2652 1572
rect 1024 34 2702 322
rect 1024 10 1618 34
<< via1 >>
rect -960 1638 -668 1914
rect -128 1666 124 1924
rect 796 1686 1048 1944
rect 1604 1702 1856 1960
rect 2376 1682 2628 1940
<< metal2 >>
rect -1084 1914 -554 2018
rect -1084 1638 -960 1914
rect -668 1638 -554 1914
rect -1084 1538 -554 1638
rect -222 1924 308 2052
rect -222 1666 -128 1924
rect 124 1666 308 1924
rect -222 1572 308 1666
rect 664 1944 1194 2062
rect 664 1686 796 1944
rect 1048 1686 1194 1944
rect 664 1582 1194 1686
rect 1548 1960 2078 2102
rect 1548 1702 1604 1960
rect 1856 1702 2078 1960
rect 1548 1622 2078 1702
rect 2310 1940 2840 2108
rect 2310 1682 2376 1940
rect 2628 1682 2840 1940
rect 2310 1628 2840 1682
use sky130_fd_pr__res_xhigh_po_0p35_K7MYC6  sky130_fd_pr__res_xhigh_po_0p35_K7MYC6_0
timestamp 1698508451
transform 1 0 27 0 1 478
box -37 -482 37 482
use sky130_fd_pr__res_xhigh_po_0p35_K7MYC6  sky130_fd_pr__res_xhigh_po_0p35_K7MYC6_1
timestamp 1698508451
transform 1 0 349 0 1 476
box -37 -482 37 482
use sky130_fd_pr__res_xhigh_po_0p35_K7MYC6  sky130_fd_pr__res_xhigh_po_0p35_K7MYC6_2
timestamp 1698508451
transform 1 0 737 0 1 476
box -37 -482 37 482
use sky130_fd_pr__res_xhigh_po_0p35_K7MYC6  sky130_fd_pr__res_xhigh_po_0p35_K7MYC6_3
timestamp 1698508451
transform 1 0 1133 0 1 472
box -37 -482 37 482
<< labels >>
rlabel metal2 -1084 1538 -960 2018 1 1
rlabel metal2 -222 1924 308 2052 1 2
rlabel metal2 664 1944 1194 2062 1 3
rlabel metal2 1548 1960 2078 2102 1 4
rlabel metal2 2310 1940 2840 2108 1 5
<< end >>

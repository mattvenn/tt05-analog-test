* divider
.lib "sky130.lib.spice" tt
.include "../lvs/netlist/tt_um_matt_divider_test.spice"

* instantiate, add VGND for VSUBS
Xcell  clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] VPWR VGND tt_um_matt_divider_test 

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* setup the transient analysis
.tran 10p 3n 0

.control
run
set color0 = white
set color1 = black
plot vgnd "uo_out[0]" "uo_out[1]" "uo_out[2]" vpwr
.endc

.end

magic
tech sky130A
magscale 1 2
timestamp 1698613918
<< via2 >>
rect 14216 19576 14556 19888
rect 15116 19640 15458 19950
rect 15952 19630 16294 19940
rect 16800 19614 17120 19986
rect 17600 19602 17996 19964
<< metal3 >>
rect 17428 21816 17492 21822
rect 15282 21752 15288 21816
rect 15352 21814 15358 21816
rect 15352 21754 17428 21814
rect 15352 21752 15358 21754
rect 17428 21746 17492 21752
rect 20208 20826 20322 20828
rect 20208 20762 20240 20826
rect 20304 20762 20322 20826
rect 16660 20078 17238 20104
rect 14986 19950 15518 20002
rect 14170 19888 14618 19934
rect 14170 19868 14216 19888
rect 14170 19570 14214 19868
rect 14556 19576 14618 19888
rect 14538 19570 14618 19576
rect 14170 19526 14618 19570
rect 14986 19572 15100 19950
rect 15458 19640 15518 19950
rect 15452 19572 15518 19640
rect 14986 19474 15518 19572
rect 15864 19966 16392 20058
rect 15864 19588 15942 19966
rect 16294 19588 16392 19966
rect 15864 19520 16392 19588
rect 16660 19582 16696 20078
rect 17198 19582 17238 20078
rect 16660 19536 17238 19582
rect 17554 19964 18048 20026
rect 17554 19602 17600 19964
rect 17996 19602 18048 19964
rect 17554 19566 18048 19602
rect 20208 17843 20322 20762
rect 20208 17779 20241 17843
rect 20305 17779 20322 17843
rect 20208 17766 20322 17779
<< via3 >>
rect 15288 21752 15352 21816
rect 17428 21752 17492 21816
rect 20240 20762 20304 20826
rect 14214 19576 14216 19868
rect 14216 19576 14538 19868
rect 14214 19570 14538 19576
rect 15100 19640 15116 19950
rect 15116 19640 15452 19950
rect 15100 19572 15452 19640
rect 15942 19940 16294 19966
rect 15942 19630 15952 19940
rect 15952 19630 16294 19940
rect 15942 19588 16294 19630
rect 16696 19986 17198 20078
rect 16696 19614 16800 19986
rect 16800 19614 17120 19986
rect 17120 19614 17198 19986
rect 16696 19582 17198 19614
rect 17600 19602 17996 19964
rect 20241 17779 20305 17843
<< metal4 >>
rect 4294 22104 4354 22304
rect 4846 22104 4906 22304
rect 5398 22104 5458 22304
rect 5950 22104 6010 22304
rect 6502 22104 6562 22304
rect 7054 22104 7114 22304
rect 7606 22104 7666 22304
rect 8158 22104 8218 22304
rect 8710 22104 8770 22304
rect 9262 22104 9322 22304
rect 9814 22104 9874 22304
rect 10366 22104 10426 22304
rect 10918 22104 10978 22304
rect 11470 22104 11530 22304
rect 12022 22104 12082 22304
rect 12574 22104 12634 22304
rect 13126 22104 13186 22304
rect 13678 22104 13738 22304
rect 14230 22104 14290 22304
rect 14782 22104 14842 22304
rect 15334 22194 15394 22304
rect 15332 22104 15394 22194
rect 15886 22146 15946 22304
rect 16438 22158 16498 22304
rect 15332 21996 15392 22104
rect 15290 21936 15392 21996
rect 15290 21817 15350 21936
rect 15287 21816 15353 21817
rect 15287 21752 15288 21816
rect 15352 21752 15353 21816
rect 15287 21751 15353 21752
rect 15120 21288 15420 21292
rect 15810 21288 15962 22146
rect 7672 20132 12790 21236
rect 15022 21138 15962 21288
rect 16376 21178 16528 22158
rect 16990 22138 17050 22304
rect 16948 21220 17100 22138
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 22104 22018 22304
rect 22510 22104 22570 22304
rect 23062 22104 23122 22304
rect 23614 22104 23674 22304
rect 24166 22104 24226 22304
rect 24718 22104 24778 22304
rect 25270 22104 25330 22304
rect 17427 21816 17493 21817
rect 17427 21752 17428 21816
rect 17492 21814 17493 21816
rect 25822 21814 25882 22304
rect 26374 22104 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 17492 21754 19108 21814
rect 20230 21754 25882 21814
rect 17492 21752 17493 21754
rect 17427 21751 17493 21752
rect 19048 21700 19108 21754
rect 20242 21620 20302 21754
rect 19050 21560 20302 21620
rect 15022 21122 15910 21138
rect 7672 19868 14692 20132
rect 15120 20016 15420 21122
rect 16184 20394 16572 21178
rect 15864 20244 16572 20394
rect 15864 20104 16396 20244
rect 16898 20150 17238 21220
rect 20242 20827 20302 21560
rect 20239 20826 20305 20827
rect 20239 20762 20240 20826
rect 20304 20762 20305 20826
rect 20239 20761 20305 20762
rect 7672 19570 14214 19868
rect 14538 19570 14692 19868
rect 7672 19274 14692 19570
rect 14986 19950 15524 20016
rect 14986 19572 15100 19950
rect 15452 19572 15524 19950
rect 15860 19966 16398 20104
rect 15860 19588 15942 19966
rect 16294 19588 16398 19966
rect 15860 19572 16398 19588
rect 16618 20078 17300 20150
rect 22610 20092 27728 21486
rect 16618 19582 16696 20078
rect 17198 19582 17300 20078
rect 14986 19484 15524 19572
rect 16618 19510 17300 19582
rect 17492 19964 27728 20092
rect 17492 19602 17600 19964
rect 17996 19602 27728 19964
rect 7672 598 12790 19274
rect 17492 18968 27728 19602
rect 20240 17843 20306 17844
rect 20240 17779 20241 17843
rect 20305 17779 20306 17843
rect 20240 17778 20306 17779
rect 20243 15172 20303 17778
rect 22610 1522 27728 18968
rect 17228 848 27728 1522
rect 17228 768 26472 848
use cap  cap_0
timestamp 1698610993
transform 1 0 13504 0 1 9908
box -318 -9140 8864 5582
use divider  divider_1
timestamp 1698571942
transform 1 0 15224 0 1 17950
box -1084 -698 2840 2108
use sky130_fd_pr__res_generic_m4_RPNQRH  sky130_fd_pr__res_generic_m4_RPNQRH_0
timestamp 1698613918
transform 1 0 19078 0 1 21665
box -30 -87 30 87
<< labels >>
flabel metal4 s 26926 22104 26986 22304 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 27478 22104 27538 22304 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 26374 22104 26434 22304 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 25270 22104 25330 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 24718 22104 24778 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 24166 22104 24226 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 23062 22104 23122 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 22510 22104 22570 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 21958 22104 22018 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 20854 22104 20914 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 20302 22104 20362 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 19750 22104 19810 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 18646 22104 18706 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 18094 22104 18154 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 17542 22104 17602 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 7606 22104 7666 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 7054 22104 7114 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 6502 22104 6562 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 5398 22104 5458 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 4846 22104 4906 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 4294 22104 4354 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 12022 22104 12082 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 11470 22104 11530 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 10918 22104 10978 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 9814 22104 9874 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 9262 22104 9322 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 8710 22104 8770 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 16438 22104 16498 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 15886 22104 15946 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 15334 22104 15394 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 14230 22104 14290 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 13678 22104 13738 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 13126 22104 13186 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal tristate
rlabel metal4 7672 598 12790 21236 1 VPWR
port 43 nsew power default
rlabel metal4 22610 848 27728 21486 1 VGND
port 44 nsew ground default
<< properties >>
string FIXED_BBOX 0 0 31464 22304
<< end >>
